/*
 * Copyright (c) 2024 Uri Shaked
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_mandelbrot_accel (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  assign uo_out  = {7'b0, o_unbounded};
  assign uio_oe  = 0;
  assign uio_out = 0;

  wire i_start = ui_in[0];
  wire [3:0] Cr_in = uio_in[3:0];
  wire [3:0] Ci_in = uio_in[7:4];

  reg o_unbounded;

  reg [31:0] Cr_next;
  reg [31:0] Ci_next;

  reg [31:0] Zr;
  reg [31:0] Zi;
  reg [31:0] Cr;
  reg [31:0] Ci;
  wire [31:0] Rr;
  wire [31:0] Ri;
  wire unbounded;

  mandelbrot_func mandelbrot (
      .Ci(Ci),
      .Cr(Cr),
      .Zr(Zr),
      .Zi(Zi),
      .Rr(Rr),
      .Ri(Ri),
      .unbounded(unbounded)
  );

  always @(posedge clk or negedge rst_n)
    if (~rst_n) begin
      Zr <= 0;
      Zi <= 0;
      Cr <= 0;
      Ci <= 0;
      Cr_next <= 0;
      Ci_next <= 0;
      o_unbounded <= 0;
    end else begin
      if (i_start) begin
        Zr <= 0;
        Zi <= 0;
        Cr <= Cr_next;
        Ci <= Ci_next;
      end else begin
        Zr <= Rr;
        Zi <= Ri;
        Cr_next <= {Cr_in, Cr_next[31:4]};
        Ci_next <= {Ci_in, Ci_next[31:4]};
        o_unbounded <= unbounded;
      end
    end

  // List all unused inputs to prevent warnings
  wire _unused = &{ena, ui_in[7:1], 1'b0};

endmodule
